//  Class: router_mcsequencer
//
class router_mcsequencer extends uvm_sequencer;
    
    `uvm_component_utils(router_mcsequencer)

    function new(string name = "router_mcsequencer", uvm_component parent = null);
      super.new(name, parent);
    endfunction
    
    
endclass: router_mcsequencer